library verilog;
use verilog.vl_types.all;
entity Top_Module_tb is
end Top_Module_tb;
