library verilog;
use verilog.vl_types.all;
entity cache_top_tb is
end cache_top_tb;
